// Benchmark "output" written by ABC on Sun Dec 24 20:15:52 2023

module output ( 
    c, d,
    F  );
  input  c, d;
  output F;
  NOR2     g0(.A(d), .B(c), .Y(F));
endmodule


