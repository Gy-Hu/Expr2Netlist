// Benchmark "output" written by ABC on Sun Dec 24 20:09:25 2023

module output ( 
    b, c,
    F  );
  input  b, c;
  output F;
  BUF_X1X1 g0(.A(b), .Y(F));
endmodule


